`timescale 1ns / 1ns
`include "alu.v"
`include "regfile.v"

module CPU(
	LEDs
	);
	
	output [7:0] LEDs;
	

endmodule
